`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/23/2023 02:54:46 PM
// Design Name: 
// Module Name: hex7seg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module hex7seg(
    input [3:0] n,
    output [6:0] s
    );
    
    m8_1 A( .in({1'b0,n[0],n[0],1'b0,1'b0,~n[0],1'b0,n[0]}), .sel(n[3:1]), .e(1'b1), .o(s[0]));
    m8_1 B( .in({1'b1,~n[0],n[0],1'b0,~n[0],n[0],1'b0,1'b0}), .sel(n[3:1]), .e(1'b1), .o(s[1]));
    m8_1 C( .in({1'b1,~n[0],1'b0,1'b0,1'b0,1'b0,~n[0],1'b0}), .sel(n[3:1]), .e(1'b1), .o(s[2]));
    m8_1 D( .in({n[0],1'b0,~n[0],n[0],n[0],~n[0],1'b0,n[0]}), .sel(n[3:1]), .e(1'b1), .o(s[3]));
    m8_1 E( .in({1'b0,1'b0,1'b0,n[0],n[0],1'b1,n[0],n[0]}), .sel(n[3:1]), .e(1'b1), .o(s[4]));
    m8_1 F( .in({1'b0,n[0],1'b0,1'b0,n[0],1'b0,1'b1,n[0]}), .sel(n[3:1]), .e(1'b1), .o(s[5]));
    m8_1 G( .in({1'b0,~n[0],1'b0,1'b0,n[0],1'b0,1'b0,1'b1}), .sel(n[3:1]), .e(1'b1), .o(s[6]));
    
//   assign s[0] = ~n[3] & ~n[2] & ~ n[1] & n[0] | ~n[3] & n[2] & ~n[1] & ~n[0] | n[3] & ~n[2] & n[1] & n[0] | n[3] & n[2] & ~n[1] & n[0];
//   assign s[1] = ~n[3] & n[2] & ~ n[1] & n[0] | ~n[3] & n[2] & n[1] & ~n[0] | n[3] & ~n[2] & n[1] & n[0] | n[3] & n[2] & ~n[1] & ~n[0] | n[3] & n[2] & n[1] & ~n[0] | n[3] & n[2] & n[1] & n[0];
//   assign s[2] = ~ n[3] & ~n[2] & n[1] & ~n[0] | n[3] & n[2] & ~n[1] & ~n[0] | n[3] & n[2] & n[1] & ~n[0] | n[3] & n[2] & n[1] & n[0];
//   assign s[3] = ~ n[3] & ~ n[2] & ~ n[1] & n[0] | ~n[3] & n[2] & ~ n[1] & ~n[0] | ~n[3] & n[2] & n[1] & n[0] | n[3] & ~n[2] & n[1] & ~n[0] | n[3] & n[2] & n[1] & n[0];
//   assign s[4] = ~ n[3] & ~n[2] & ~n[1] & n[0] | ~n[3] & ~n[2] & n[1] & n[0] | ~n[3] & n[2] & ~n[1] & ~n[0] | ~n[3] & n[2] & ~n[1] & n[0] | ~n[3] & n[2] & n[1] & n[0] | n[3] & ~n[2] & ~n[1] & n[0];
//   assign s[5] = ~n[3] & ~n[2] & ~n[1] & n[0] | ~n[3] & ~n[2] & n[1] & ~n[0] | ~n[3] & ~n[2] & n[1] & n[0] | ~n[3] & n[2] & n[1] & n[0] | n[3] & n[2] & ~n[1] & n[0]; 
//   assign s[6] = ~n[3] & ~n[2] & ~n[1] & ~n[0] | ~n[3] & ~n[2] & ~n[1] & n[0] | ~n[3] & n[2] & n[1] & n[0] |n[3] & n[2] & ~n[1] & ~n[0];
endmodule
